`define SYS_CLK 50_000_000

module top_module (
    input start,
    input skip,
    input reset,
    input clk,
    input [2:0] weight,
    input [1:0] calories,
    input [1:0] MET,
    input gender,
    output [4:0] seg_sel,
    output [7:0] seg_data,
    output buzzer_out
    );

    wire [1:0] state_w;
    wire [5:0] timer_w;
    wire [7:0] curr_idx_w;
    wire act_buz_w;
    wire buz_mode_w;
    wire [8:0] total_workouts;
    wire [7:0] total_workouts_8bit;
    
    combinational_circuit calc1(
        .input_bits({weight, calories, MET, gender}),
        .T3(total_workouts_8bit)
    );
    assign total_workouts = {1'b0, total_workouts_8bit};

    workout_fsm f1(
        .start_btn(start),
        .skip_btn(skip),
        .reset_btn(reset),
        .clk(clk),
        .total_count_in(total_workouts),
        .state(state_w),
        .timer(timer_w),
        .curr_idx(curr_idx_w),
        .buz_pulse(act_buz_w),
        .buz_mode(buz_mode_w)
    );

    wire short_beep, long_beep;
    assign short_beep = act_buz_w & ~buz_mode_w;
    assign long_beep = act_buz_w & buz_mode_w;
    
    BuzzerControllerParamR b1(
        .clk(clk),
        .rst(~reset),
        .shortBeepTrig(short_beep),
        .longBeepTrig(long_beep),
        .buzzer(buzzer_out)
    );

    wire [8:0] to_show;
    assign to_show = (state_w == 2'b00) ? total_workouts : {1'b0, curr_idx_w};

    //---------- New 7-Segment Display Logic Wires ----------
    wire [3:0] timer_tens, timer_ones;   //BCD
    wire [3:0] workout_tens, workout_ones;  //BCD
    wire [3:0] selected_digit;
    wire [2:0] refresh_counter_wire;
    wire refresh_clk;

    //---------- Clock Divider for Display Refresh (~760 Hz) ----------
    reg [15:0] refresh_clk_counter = 0;
    assign refresh_clk = refresh_clk_counter[15];  // clock output
    always @(posedge clk) begin
        refresh_clk_counter <= refresh_clk_counter + 1;
    end

    //---------- New Module Instantiations for Display ----------
    refreshCounter rc_inst (
        .refresh_clock(refresh_clk),
        .refreshCounter(refresh_counter_wire)
    );

    digit_multiplexer dm_inst (
        .refreshCounter(refresh_counter_wire),
        .SEG_SEL(seg_sel)
    );
    
    bin_to_bcd timer_converter (
        .binary(timer_w), // timer is 6-bit, fits in 8-bit input
        .tens(timer_tens),
        .ones(timer_ones)
    );

    bin_to_bcd workout_converter (
        .binary(to_show[7:0]),
        .tens(workout_tens),
        .ones(workout_ones)
    );

    BCDcontrol bcd_ctrl_inst (
        .digit1(workout_ones),
        .digit2(workout_tens),
        .digit3(timer_ones),
        .digit4(timer_tens),
        .refreshCounter(refresh_counter_wire),
        .one_digit(selected_digit)
    );
    
    bcd2seven_seg seg_decoder_inst (
        .digit(selected_digit),
        .SEG_DATA(seg_data)
    );

endmodule




module combinational_circuit (
    input  [7:0] input_bits,
    output [7:0] T3
    );

    wire w2 = input_bits[7];
    wire w1 = input_bits[6];
    wire w0 = input_bits[5];
    wire c1 = input_bits[4];
    wire c0 = input_bits[3];
    wire M1 = input_bits[2];
    wire M0 = input_bits[1];
    wire G  = input_bits[0];

    wire [7:0] T1;

    assign T1[0] = (~w2 & ~c1 & c0 & w1 & w0) | (c1 & c0 & w1 & ~w0) | (~w2 & ~c0 & w1 & ~w0) | (w2 & c0 & ~w0) | (w2 & ~c1 & ~w0) | (w2 & ~c0 & w1 & w0);
    assign T1[1] = (~w2 & c0 & w1) | (~w2 & ~c1 & w1) | (~c1 & c0 & w1) | (~c0 & ~w1 & w0) | (w2 & ~c1 & c0 & ~w0) | (w2 & c1 & ~c0 & w1) | (w2 & ~c0 & w1 & ~w0);
    assign T1[2] = (~c1 & c0 & ~w1 & w0) | (c1 & c0 & w1 & w0) | (~c1 & c0 & w1 & ~w0) | (~w2 & c1 & ~c0 & ~w1 ) | (~w2 & ~c0 & ~w1 & ~w0) | (~w2 & ~c1 & ~c0 & w1 & w0) | (w2 & c1 & ~w1 & ~w0) | (w2 & c0 & w1 & ~w0) | (w2 & ~c1 & ~w1 & w0);
    assign T1[3] = (w2 & ~w1 & w0 ) | (w2 & ~c0 & w1 & w0 ) | (c1 & c0 & ~w1 & w0) | (c1 & c0 & w1 & ~w0) | (~c1 & ~c0 & w1 & ~w0) | (~w2 & ~c1 & c0 & w1 & w0) | (~w2 & ~c1 & ~w1 & ~w0);
    assign T1[4] = (~c0 & ~w2 & ~w1) | (~w2 & ~w1 & ~w0) | (~c1 & c0 & w1 & ~w0) | (~c0 & w2 & w1 & ~w0 ) | (c1 & ~w2 & w1 & w0 ) | (~c1 & w2 & w0) | (w2 & ~w1 & w0);
    assign T1[5] = (~c1 & ~c0 & ~w2) | (~w2 & ~w1 & ~w0) | (~c1 & ~w2 & ~w1 ) | (c1 & c0 & ~w2 & ~w0 ) | (c0 & w2 & w1) | (~c0 & w2 & ~w1 & ~w0) | (~c0 & ~w2 & w1 & w0) | (c0 & w2 & w0);
    assign T1[6] = (~c1 & c0 & ~w2) | (~c1 & c0 & ~w1 & ~w0) | (c0 & ~w2 & ~w1) | (c1 & w2 & w1) | (c1 & w2 & w0) | (c1 & ~c0 & w2) | (c1 & ~c0 & w1 & w0);
    assign T1[7] = (c1 & c0 & ~w2) | (c1 & ~w2 & ~w0)  | (c1 & ~w2 & ~w1) | (c1 & c0 & ~w1 & ~w0);

    wire [7:0] T1_shifted = {3'b000, T1[7:3]};
    wire [7:0] T1_woman;
    wire [8:0] carry;
    assign carry[0] = 0;

    full_adder fa0 (.a(T1[0]), .b(T1_shifted[0]), .cin(carry[0]), .sum(T1_woman[0]), .cout(carry[1]));
    full_adder fa1 (.a(T1[1]), .b(T1_shifted[1]), .cin(carry[1]), .sum(T1_woman[1]), .cout(carry[2]));
    full_adder fa2 (.a(T1[2]), .b(T1_shifted[2]), .cin(carry[2]), .sum(T1_woman[2]), .cout(carry[3]));
    full_adder fa3 (.a(T1[3]), .b(T1_shifted[3]), .cin(carry[3]), .sum(T1_woman[3]), .cout(carry[4]));
    full_adder fa4 (.a(T1[4]), .b(T1_shifted[4]), .cin(carry[4]), .sum(T1_woman[4]), .cout(carry[5]));
    full_adder fa5 (.a(T1[5]), .b(T1_shifted[5]), .cin(carry[5]), .sum(T1_woman[5]), .cout(carry[6]));
    full_adder fa6 (.a(T1[6]), .b(T1_shifted[6]), .cin(carry[6]), .sum(T1_woman[6]), .cout(carry[7]));
    full_adder fa7 (.a(T1[7]), .b(T1_shifted[7]), .cin(carry[7]), .sum(T1_woman[7]), .cout(carry[8]));

    wire [7:0] T2;
    assign T2[0] = (~G & T1[0]) | (G & T1_woman[0]);
    assign T2[1] = (~G & T1[1]) | (G & T1_woman[1]);
    assign T2[2] = (~G & T1[2]) | (G & T1_woman[2]);
    assign T2[3] = (~G & T1[3]) | (G & T1_woman[3]);
    assign T2[4] = (~G & T1[4]) | (G & T1_woman[4]);
    assign T2[5] = (~G & T1[5]) | (G & T1_woman[5]);
    assign T2[6] = (~G & T1[6]) | (G & T1_woman[6]);
    assign T2[7] = (~G & T1[7]) | (G & T1_woman[7]);

    wire [7:0] shift0 = T2;
    wire [7:0] shift1 = {1'b0, T2[7:1]};
    wire [7:0] shift2 = {2'b00, T2[7:2]};
    wire [7:0] shift3 = {3'b000, T2[7:3]};

    mux4x1 mux0 (.in0(shift0[0]), .in1(shift1[0]), .in2(shift2[0]), .in3(shift3[0]), .sel({M1, M0}), .out(T3[0]));
    mux4x1 mux1 (.in0(shift0[1]), .in1(shift1[1]), .in2(shift2[1]), .in3(shift3[1]), .sel({M1, M0}), .out(T3[1]));
    mux4x1 mux2 (.in0(shift0[2]), .in1(shift1[2]), .in2(shift2[2]), .in3(shift3[2]), .sel({M1, M0}), .out(T3[2]));
    mux4x1 mux3 (.in0(shift0[3]), .in1(shift1[3]), .in2(shift2[3]), .in3(shift3[3]), .sel({M1, M0}), .out(T3[3]));
    mux4x1 mux4 (.in0(shift0[4]), .in1(shift1[4]), .in2(shift2[4]), .in3(shift3[4]), .sel({M1, M0}), .out(T3[4]));
    mux4x1 mux5 (.in0(shift0[5]), .in1(shift1[5]), .in2(shift2[5]), .in3(shift3[5]), .sel({M1, M0}), .out(T3[5]));
    mux4x1 mux6 (.in0(shift0[6]), .in1(shift1[6]), .in2(shift2[6]), .in3(shift3[6]), .sel({M1, M0}), .out(T3[6]));
    mux4x1 mux7 (.in0(shift0[7]), .in1(shift1[7]), .in2(shift2[7]), .in3(shift3[7]), .sel({M1, M0}), .out(T3[7]));

endmodule


module full_adder (
    input a, b, cin,
    output sum, cout
);
    assign sum  = a ^ b ^ cin;
    assign cout = (a & b) | (a & cin) | (b & cin);
endmodule


module mux4x1 (
    input in0, in1, in2, in3,
    input [1:0] sel,
    output out
    );
    wire n0, n1, s0, s1, s2, s3;
    not (n0, sel[0]);
    not (n1, sel[1]);
    and (s0, n1, n0, in0);
    and (s1, n1, sel[0], in1);
    and (s2, sel[1], n0, in2);
    and (s3, sel[1], sel[0], in3);
    or  (out, s0, s1, s2, s3);
endmodule


module clk_en_gen #(parameter DIVIDER = `SYS_CLK)(
    input clk,
    input reset_n,
    output reg clk_en
    );
    reg [31:0] ctr;
    always @(posedge clk or negedge reset_n) begin
        if (~reset_n) begin
            ctr <= 0;
            clk_en <= 0;
        end else begin
            if (ctr == DIVIDER - 1) begin
                ctr <= 0;
                clk_en <= 1;
            end else begin
                ctr <= ctr + 1;
                clk_en <= 0;
            end
        end
    end
endmodule


module debouncer(
    input clk,
    input rst, 
    input noisy_btn,
    output reg clean_btn
    );
    
    reg bit0;
    reg bit1;
    
    always@(posedge clk or posedge rst) begin
        if(rst) begin
            bit0 <= 1'b1;
            bit1 <= 1'b1;
            clean_btn <= 1'b1;
        end else begin
            bit0 <= noisy_btn;
            bit1 <= bit0;
            clean_btn <= bit1 & bit0;
        end
    end
endmodule



module ButtonCond #(parameter ACTIVE_LOW=1)(
    input  clk,
    input rst,
    input btn_in,
    output reg press
    );
    wire lvl_raw;
    debouncer udb (
        .clk(clk), 
        .rst(rst), 
        .noisy_btn(btn_in), 
        .clean_btn(lvl_raw)
    );
    wire lvl_norm = ACTIVE_LOW ? ~lvl_raw : lvl_raw;
    reg  prev;
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            prev<=1'b0;
            press<=1'b0;
        end else begin
            press <= (lvl_norm & ~prev);
            prev <= lvl_norm;
        end
    end
endmodule


module fsm_core_logic(
    input clk,
    input reset_n,
    input start_edge,
    input skip_edge,
    input reset_edge,
    input clk_en_rising,
    input [8:0] total_count_in,
    output reg [1:0] state = 2'b00,
    output reg [5:0] timer = 6'b101101,
    output reg [7:0] curr_idx = 0,
    output reg buz_pulse = 1'b0,
    output reg buz_mode = 0
    );
    localparam IDLE = 2'b00, EXERCISE = 2'b01, REST = 2'b10;
    
    always @(posedge clk or negedge reset_n) begin
        if (~reset_n) begin
            state        <= IDLE;
            timer        <= 6'b101101;
            curr_idx     <= 0;
            buz_pulse    <= 1'b1;
            buz_mode     <= 1'b0;
        end else begin
            buz_pulse <= 1'b0;
            if (reset_edge) begin // Global reset condition
                state <= IDLE;
                curr_idx <= 0;
            end else begin
                case (state)
                    IDLE: begin
                        timer        <= 6'b101101;
                        if (start_edge && total_count_in > 0) begin
                            curr_idx     <= total_count_in; 
                            state        <= EXERCISE;
                        end
                    end
                    EXERCISE: begin
                        if (skip_edge) begin
                            if (curr_idx > 1)
                                curr_idx <= curr_idx - 1;
                            else
                                state <= IDLE;
                            timer     <= 6'b101101;
                            buz_pulse <= 1'b1;
                        end else if (clk_en_rising) begin
                            if (timer == 1) begin
                                state     <= REST;
                                timer     <= 6'b001111;
                                buz_pulse <= 1'b1;
                            end else if (timer != 0) begin
                                timer <= timer - 1;
                            end 
                        end
                    end
                    REST: begin
                        if (skip_edge) begin
                            if (curr_idx > 1)
                                curr_idx <= curr_idx - 1;
                            else
                                state <= IDLE;
                            state     <= EXERCISE;
                            timer     <= 6'b101101;
                            buz_pulse <= 1'b1;
                        end else if (clk_en_rising) begin
                            if (timer == 1) begin
                                if (curr_idx <= 1) begin // This was the last workout
                                    state     <= IDLE;
                                    curr_idx  <= 0;
                                    buz_pulse <= 1'b1;
                                    buz_mode  <= 1'b1;
                                end else begin
                                    curr_idx  <= curr_idx - 1; 
                                    state     <= EXERCISE;
                                    timer     <= 6'b101101;
                                    buz_pulse <= 1'b1;
                                end
                            end else if (timer != 0) begin
                                timer <= timer - 1;
                            end
                        end
                    end
                endcase
            end
        end
    end
endmodule


module workout_fsm(
    input start_btn,
    input skip_btn,
    input reset_btn,
    input clk,
    input [8:0] total_count_in,
    output [1:0] state,
    output [5:0] timer,
    output [7:0] curr_idx,
    output buz_pulse,
    output buz_mode
    );
    wire start_edge, skip_edge, reset_edge;
    wire clk_out;

    ButtonCond #(.ACTIVE_LOW(1'b1))
      bc_start (.clk(clk), .rst(~reset_btn), .btn_in(start_btn), .press(start_edge));
    ButtonCond #(.ACTIVE_LOW(1'b1))
      bc_skip  (.clk(clk), .rst(~reset_btn), .btn_in(skip_btn),  .press(skip_edge));
    ButtonCond #(.ACTIVE_LOW(1'b1))
      bc_reset (.clk(clk), .rst(~reset_btn), .btn_in(reset_btn), .press(reset_edge));
    
    clk_en_gen #(.DIVIDER(`SYS_CLK)) clkgen (
        .clk(clk),
        .reset_n(reset_btn),
        .clk_en(clk_out)
    );
    
    fsm_core_logic fcl (
        .clk(clk),
        .reset_n(reset_btn),
        .start_edge(start_edge),
        .skip_edge(skip_edge),
        .reset_edge(reset_edge),
        .clk_en_rising(clk_out),
        .total_count_in(total_count_in),
        .state(state),
        .timer(timer),
        .curr_idx(curr_idx),
        .buz_pulse(buz_pulse),
        .buz_mode(buz_mode)
    );
endmodule


module BuzzerControllerParamR(
    input clk,
    input rst,
    input shortBeepTrig,
    input longBeepTrig,
    output buzzer
    );
    localparam [25:0] SHORT_CYC=26'd10000000;  // ~0.20 s
    localparam [25:0] LONG_CYC =26'd30000000; // ~0.60 s
    localparam [15:0] SHORT_DIV=16'd24999;   // ~1 kHz
    localparam [15:0] LONG_DIV =16'd12499;    // ~2 kHz
    
    reg buzzReq; reg [25:0] cntDur;
    reg [15:0] divCnt, divSel;
    reg sq;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            buzzReq<=0;
            cntDur<=0;
            divCnt<=0;
            divSel<=SHORT_DIV;
            sq<=0;
        end else begin
            if (longBeepTrig) begin
                buzzReq<=1;
                cntDur<=LONG_CYC;
                divSel<=LONG_DIV;
            end else if (shortBeepTrig) begin
                buzzReq<=1;
                cntDur<=SHORT_CYC;
                divSel<=SHORT_DIV;
            end else if (cntDur!=0) begin
                cntDur<=cntDur-1;
                buzzReq<=1;
            end else begin
                buzzReq<=0;
            end
            if (!buzzReq) begin
                divCnt<=0;
                sq<=0;
            end else if (divCnt==divSel) begin
                divCnt<=0;
                sq<=~sq;
            end else
                divCnt<=divCnt+1;
        end
    end
    assign buzzer = sq;
endmodule

//---------- New Display Modules ----------


module bcd2seven_seg ( 
    input [3:0] digit, 
    output reg [7:0] SEG_DATA = 0
); 
    always @(digit)
    begin 
        case(digit) 
            4'd0: SEG_DATA = 8'b00111111; 
            4'd1: SEG_DATA = 8'b00000110; 
            4'd2: SEG_DATA = 8'b01011011;
            4'd3: SEG_DATA = 8'b01001111; 
            4'd4: SEG_DATA = 8'b01100110; 
            4'd5: SEG_DATA = 8'b01101101; 
            4'd6: SEG_DATA = 8'b01111101; 
            4'd7: SEG_DATA = 8'b00000111; 
            4'd8: SEG_DATA = 8'b01111111;
            4'd9: SEG_DATA = 8'b01101111; 
            default: SEG_DATA = 8'b00000000; // Invalid input (all segments off)
        endcase 
    end 
endmodule 



module BCDcontrol (
    input [3:0] digit1,  // rightmost digit
    input [3:0] digit2,
    input [3:0] digit3,
    input [3:0] digit4,  // leftmost digit
    input [2:0] refreshCounter,
    output reg [3:0] one_digit = 0  // digit to be displayed
);
    always @(refreshCounter) begin
        case (refreshCounter)
            2'd0: one_digit = digit1;
            2'd1: one_digit = digit2;
            2'd2: one_digit = digit3;
            2'd3: one_digit = digit4;
            default: one_digit = digit1;
        endcase
    end
endmodule



module refreshCounter (
    input refresh_clock,
    output reg [2:0] refreshCounter = 0
);
    always @(posedge refresh_clock) begin
        if(refreshCounter == 3'b101)
            refreshCounter <= 3'b000;
        else
            refreshCounter <= refreshCounter + 1;
    end
endmodule


module digit_multiplexer (
    input [2:0] refreshCounter,
    output reg [4:0] SEG_SEL = 0
);
    always @(refreshCounter) begin
        case (refreshCounter)
            2'd0: SEG_SEL = 5'b00010; // activate rightmost digit
            2'd1: SEG_SEL = 5'b00100;
            2'd2: SEG_SEL = 5'b01000;
            2'd3: SEG_SEL = 5'b00001; // activate leftmost digit
            default: SEG_SEL = 5'b00000;
        endcase
    end
endmodule

module bin_to_bcd (
    input [7:0] binary,
    output reg [3:0] tens,
    output reg [3:0] ones
);
    integer i;
    reg [7:0] bcd;   
    always @(*) begin 
        bcd = 0;
        for (i = 0; i < 8; i = i + 1) begin
            if (bcd[3:0] >= 5)
                bcd[3:0] = bcd[3:0] + 3;
            if (bcd[7:4] >= 5)
                bcd[7:4] = bcd[7:4] + 3;
            bcd = {bcd[6:0], binary[7-i]};
        end
        tens = bcd[7:4];
        ones = bcd[3:0];
    end
endmodule